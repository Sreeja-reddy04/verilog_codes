module full_adder(a_in,
                  b_in,
		  c_in,
		  sum_out,
		  carry_out);

   //Step1 : Write down the directions for the ports	      

   //Step2 : Declare the internal wires    

   //Step3 : Instantiate the Half-Adders using name-based port mapping			 

   //Step4 : Instantiate the OR gate


endmodule

