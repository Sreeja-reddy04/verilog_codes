`timescale 1ns / 1ps

module jkff_tb;

	// Inputs
	reg j;
	reg k;
	reg clk;
	reg rst;

	// Outputs
	wire q;
	wire qb;
	integer a,b;

	// Instantiate the Unit Under Test (UUT)
	jff uut (
		.j(j), 
		.k(k), 
		.clk(clk), 
		.rst(rst), 
		.q(q), 
		.qb(qb)
	);
	
	always
	begin
	#5 clk = ('b0);
	#5 clk = ~clk;
	end
	
	task r();
	begin
	@(negedge clk);
	rst = 1'b1;
	@(negedge clk);
	rst = 1'b0;
	end
	endtask
	
	task in(input a,b);
	begin
	j=a;
	k=b;
	end
	endtask
	
	initial
	begin
	r;
	in(1'b1,1'b0);
	in(1'b0,1'b1);
	in(1'b0,1'b0);
	in(1'b1,1'b1);
	
	
	//initial begin
		// Initialize Inputs
		/*j = 0;
		k = 0;
		clk = 0;
		rst = 0;*/

		// Wait 100 ns for global reset to finish
		//#100;
        
		// Add stimulus here

	end
      
endmodule

